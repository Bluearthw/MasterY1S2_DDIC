/esat/micas-data/data/design/generic/Cadence_kits_2023/GPDK045/gsclib045_all_v4.7/gsclib045_lvt/lef/gsclib045_lvt_macro.lef